import uvm_pkg::*;

class A extends uvm_component;
	function new(string name);
		super.new(name, null);
	endfunction

	task run_phase(uvm_phase phase);
		$display("A::run_phase HELLO A.");
	endtask
endclass

class B extends uvm_component;
	function new(string name);
		super.new(name, null);
	endfunction

	task run_phase(uvm_phase phase);
		$display("B::run_phase HELLO B.");
	endtask
endclass

// C will not be phased because it is not contained in uvm_top
class C extends uvm_component;
	function new(string name);
		super.new(name, null);
	endfunction

	task run_phase(uvm_phase phase);
		$display("C::run_phase HELLO C.");
	endtask
endclass

module test;
	A a;
	B b;

	initial 
	begin
		a = new("uA");
		b = new("uB");
		run_test();
	end
endmodule

