module top;
	initial 
		$hello();
endmodule

